-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Saturday, April 04, 2015 12:21:38 �й���׼ʱ��

